library ieee; 
use ieee.std_logic_1164.all; 
use work.components.all;  

entity FSM_Controller is 
	port(		: in std_logic;
				: out std_logic);
end FSM_Controller;


ARCHITECTURE struc_behavior OF FSM_Controller is
BEGIN

--- 2to1Mux ---


--- bitwise_and ---


end struc_behavior;